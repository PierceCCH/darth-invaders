`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:58:41 03/08/2023 
// Design Name: 
// Module Name:    components 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module components(
    input d_left,
    input d_right,
    input d_fire,
    input d_reset,
    output proj_xcoord,
    output proj_ycoord,
    output ship_xcoord,
    output ship_ycoord
    );


endmodule
